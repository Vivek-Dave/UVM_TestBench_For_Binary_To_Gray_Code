class bintogray_sequencer extends uvm_sequencer#(bintogray_sequence_item);
  //----------------------------------------------------------------------------
  `uvm_component_utils(bintogray_sequencer)  
  //----------------------------------------------------------------------------

  //----------------------------------------------------------------------------
  function new(string name="bintogray_sequencer",uvm_component parent);  
    super.new(name,parent);
  endfunction
  //----------------------------------------------------------------------------
  
endclass:bintogray_sequencer

