
interface intf();
    // ------------------- port declaration-------------------------------------
    logic [7:0]  in;
    logic [7:0] out;
    //--------------------------------------------------------------------------
endinterface

